// Dummy user_defines.v for demo
module user_defines();
endmodule 